library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity de2-cpu is
	port(		: in --type
	;
				: out --type
	);
end de2-cpu;